-- Copyright (C) 2022  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 22.1std.0 Build 915 10/25/2022 SC Lite Edition"
-- CREATED		"Mon Jan 13 20:30:24 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY zegarek IS 
	PORT
	(
		S :  IN  STD_LOGIC;
		U :  IN  STD_LOGIC;
		CLK_50MHz :  IN  STD_LOGIC;
		s_sekunda :  IN  STD_LOGIC;
		clr :  IN  STD_LOGIC;
		pin_name1 :  OUT  STD_LOGIC;
		Seg_out0 :  OUT  STD_LOGIC;
		Seg_out1 :  OUT  STD_LOGIC;
		Seg_out2 :  OUT  STD_LOGIC;
		Seg_out3 :  OUT  STD_LOGIC;
		Seg_out4 :  OUT  STD_LOGIC;
		Seg_out5 :  OUT  STD_LOGIC;
		Seg_out6 :  OUT  STD_LOGIC;
		Seg_out10 :  OUT  STD_LOGIC;
		Seg_out11 :  OUT  STD_LOGIC;
		Seg_out12 :  OUT  STD_LOGIC;
		Seg_out13 :  OUT  STD_LOGIC;
		Seg_out14 :  OUT  STD_LOGIC;
		Seg_out15 :  OUT  STD_LOGIC;
		Seg_out16 :  OUT  STD_LOGIC;
		Seg_out20 :  OUT  STD_LOGIC;
		Seg_out21 :  OUT  STD_LOGIC;
		Seg_out22 :  OUT  STD_LOGIC;
		Seg_out23 :  OUT  STD_LOGIC;
		Seg_out24 :  OUT  STD_LOGIC;
		Seg_out25 :  OUT  STD_LOGIC;
		Seg_out26 :  OUT  STD_LOGIC;
		Seg_out30 :  OUT  STD_LOGIC;
		Seg_out31 :  OUT  STD_LOGIC;
		Seg_out32 :  OUT  STD_LOGIC;
		Seg_out33 :  OUT  STD_LOGIC;
		Seg_out34 :  OUT  STD_LOGIC;
		Seg_out35 :  OUT  STD_LOGIC;
		Seg_out36 :  OUT  STD_LOGIC
	);
END zegarek;

ARCHITECTURE bdf_type OF zegarek IS 

COMPONENT edgeing
	PORT(clk : IN STD_LOGIC;
		 D_in : IN STD_LOGIC;
		 Q : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT preskalervhdl
	PORT(CLK_50MHz : IN STD_LOGIC;
		 CLK_10Hz : OUT STD_LOGIC;
		 CLK_1Hz : OUT STD_LOGIC;
		 CLK_1_60Hz : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT liczniktrzy
	PORT(CLK_50MHz : IN STD_LOGIC;
		 CLK_1Hz : IN STD_LOGIC;
		 U : IN STD_LOGIC;
		 OUTPUT : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT licznik_10
	PORT(clk : IN STD_LOGIC;
		 en : IN STD_LOGIC;
		 clr : IN STD_LOGIC;
		 rco : OUT STD_LOGIC;
		 Q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT bcd_to_7seg
	PORT(BCD_in : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Seg_out : OUT STD_LOGIC_VECTOR(0 TO 6)
	);
END COMPONENT;

SIGNAL	Q0 :  STD_LOGIC;
SIGNAL	Q1 :  STD_LOGIC;
SIGNAL	Q10 :  STD_LOGIC;
SIGNAL	Q11 :  STD_LOGIC;
SIGNAL	Q12 :  STD_LOGIC;
SIGNAL	Q13 :  STD_LOGIC;
SIGNAL	Q2 :  STD_LOGIC;
SIGNAL	Q20 :  STD_LOGIC;
SIGNAL	Q21 :  STD_LOGIC;
SIGNAL	Q22 :  STD_LOGIC;
SIGNAL	Q23 :  STD_LOGIC;
SIGNAL	Q3 :  STD_LOGIC;
SIGNAL	Q30 :  STD_LOGIC;
SIGNAL	Q31 :  STD_LOGIC;
SIGNAL	Q32 :  STD_LOGIC;
SIGNAL	Q33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	TFF_inst321 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	TFF_inst322 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC_VECTOR(0 TO 6);
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC_VECTOR(0 TO 6);
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC_VECTOR(0 TO 6);
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC_VECTOR(0 TO 6);

SIGNAL	GDFX_TEMP_SIGNAL_3 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_7 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_2 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_6 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_5 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_4 :  STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN 
Seg_out0 <= SYNTHESIZED_WIRE_60(0);
Seg_out1 <= SYNTHESIZED_WIRE_60(1);
Seg_out2 <= SYNTHESIZED_WIRE_60(2);
Seg_out3 <= SYNTHESIZED_WIRE_60(3);
Seg_out4 <= SYNTHESIZED_WIRE_60(4);
Seg_out5 <= SYNTHESIZED_WIRE_60(5);
Seg_out6 <= SYNTHESIZED_WIRE_60(6);
Seg_out10 <= SYNTHESIZED_WIRE_61(0);
Seg_out11 <= SYNTHESIZED_WIRE_61(1);
Seg_out12 <= SYNTHESIZED_WIRE_61(2);
Seg_out13 <= SYNTHESIZED_WIRE_61(3);
Seg_out14 <= SYNTHESIZED_WIRE_61(4);
Seg_out15 <= SYNTHESIZED_WIRE_61(5);
Seg_out16 <= SYNTHESIZED_WIRE_61(6);
Seg_out20 <= SYNTHESIZED_WIRE_62(0);
Seg_out21 <= SYNTHESIZED_WIRE_62(1);
Seg_out22 <= SYNTHESIZED_WIRE_62(2);
Seg_out23 <= SYNTHESIZED_WIRE_62(3);
Seg_out24 <= SYNTHESIZED_WIRE_62(4);
Seg_out25 <= SYNTHESIZED_WIRE_62(5);
Seg_out26 <= SYNTHESIZED_WIRE_62(6);
Seg_out30 <= SYNTHESIZED_WIRE_63(0);
Seg_out31 <= SYNTHESIZED_WIRE_63(1);
Seg_out32 <= SYNTHESIZED_WIRE_63(2);
Seg_out33 <= SYNTHESIZED_WIRE_63(3);
Seg_out34 <= SYNTHESIZED_WIRE_63(4);
Seg_out35 <= SYNTHESIZED_WIRE_63(5);
Seg_out36 <= SYNTHESIZED_WIRE_63(6);

Q33 <= GDFX_TEMP_SIGNAL_3(3);
Q32 <= GDFX_TEMP_SIGNAL_3(2);
Q31 <= GDFX_TEMP_SIGNAL_3(1);
Q30 <= GDFX_TEMP_SIGNAL_3(0);

GDFX_TEMP_SIGNAL_7 <= (Q33 & Q32 & Q31 & Q30);
Q23 <= GDFX_TEMP_SIGNAL_2(3);
Q22 <= GDFX_TEMP_SIGNAL_2(2);
Q21 <= GDFX_TEMP_SIGNAL_2(1);
Q20 <= GDFX_TEMP_SIGNAL_2(0);

GDFX_TEMP_SIGNAL_6 <= (Q23 & Q22 & Q21 & Q20);
Q13 <= GDFX_TEMP_SIGNAL_1(3);
Q12 <= GDFX_TEMP_SIGNAL_1(2);
Q11 <= GDFX_TEMP_SIGNAL_1(1);
Q10 <= GDFX_TEMP_SIGNAL_1(0);

GDFX_TEMP_SIGNAL_5 <= (Q13 & Q12 & Q11 & Q10);
Q3 <= GDFX_TEMP_SIGNAL_0(3);
Q2 <= GDFX_TEMP_SIGNAL_0(2);
Q1 <= GDFX_TEMP_SIGNAL_0(1);
Q0 <= GDFX_TEMP_SIGNAL_0(0);

GDFX_TEMP_SIGNAL_4 <= (Q3 & Q2 & Q1 & Q0);


b2v_inst : edgeing
PORT MAP(clk => CLK_50MHz,
		 D_in => SYNTHESIZED_WIRE_0,
		 Q => SYNTHESIZED_WIRE_57);


SYNTHESIZED_WIRE_6 <= CLK_50MHz AND SYNTHESIZED_WIRE_1;


b2v_inst12 : preskalervhdl
PORT MAP(CLK_50MHz => CLK_50MHz,
		 CLK_1Hz => SYNTHESIZED_WIRE_55);


SYNTHESIZED_WIRE_8 <= TFF_inst321 AND SYNTHESIZED_WIRE_54;


SYNTHESIZED_WIRE_58 <= Q11 AND Q12;


b2v_inst18 : liczniktrzy
PORT MAP(CLK_50MHz => CLK_50MHz,
		 CLK_1Hz => SYNTHESIZED_WIRE_55,
		 U => SYNTHESIZED_WIRE_56,
		 OUTPUT => SYNTHESIZED_WIRE_1);


SYNTHESIZED_WIRE_56 <= NOT(U);



PROCESS(CLK_50MHz)
VARIABLE pin_name1_synthesized_var : STD_LOGIC;
BEGIN
IF (RISING_EDGE(CLK_50MHz)) THEN
	pin_name1_synthesized_var := pin_name1_synthesized_var XOR SYNTHESIZED_WIRE_54;
END IF;
	pin_name1 <= pin_name1_synthesized_var;
END PROCESS;


b2v_inst21 : preskalervhdl
PORT MAP(CLK_50MHz => SYNTHESIZED_WIRE_6,
		 CLK_10Hz => SYNTHESIZED_WIRE_7);


b2v_inst22 : preskalervhdl
PORT MAP(CLK_50MHz => CLK_50MHz,
		 CLK_1_60Hz => SYNTHESIZED_WIRE_54);


SYNTHESIZED_WIRE_29 <= NOT(s_sekunda);



SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_9 <= SYNTHESIZED_WIRE_55 AND TFF_inst322;


b2v_inst29 : licznik_10
PORT MAP(clk => CLK_50MHz,
		 en => SYNTHESIZED_WIRE_12,
		 clr => SYNTHESIZED_WIRE_57,
		 rco => SYNTHESIZED_WIRE_14,
		 Q => GDFX_TEMP_SIGNAL_0);


SYNTHESIZED_WIRE_27 <= NOT(S);



b2v_inst30 : licznik_10
PORT MAP(clk => CLK_50MHz,
		 en => SYNTHESIZED_WIRE_14,
		 clr => SYNTHESIZED_WIRE_15,
		 Q => GDFX_TEMP_SIGNAL_1);


SYNTHESIZED_WIRE_0 <= NOT(clr);



b2v_inst32 : licznik_10
PORT MAP(clk => CLK_50MHz,
		 en => SYNTHESIZED_WIRE_58,
		 clr => SYNTHESIZED_WIRE_59,
		 rco => SYNTHESIZED_WIRE_24,
		 Q => GDFX_TEMP_SIGNAL_2);


PROCESS(CLK_50MHz)
VARIABLE TFF_inst321_synthesized_var : STD_LOGIC;
BEGIN
IF (RISING_EDGE(CLK_50MHz)) THEN
	TFF_inst321_synthesized_var := TFF_inst321_synthesized_var XOR SYNTHESIZED_WIRE_18;
END IF;
	TFF_inst321 <= TFF_inst321_synthesized_var;
END PROCESS;


PROCESS(CLK_50MHz)
VARIABLE TFF_inst322_synthesized_var : STD_LOGIC;
BEGIN
IF (RISING_EDGE(CLK_50MHz)) THEN
	TFF_inst322_synthesized_var := TFF_inst322_synthesized_var XOR SYNTHESIZED_WIRE_19;
END IF;
	TFF_inst322 <= TFF_inst322_synthesized_var;
END PROCESS;


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_58;


SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_23;


b2v_inst35 : licznik_10
PORT MAP(clk => CLK_50MHz,
		 en => SYNTHESIZED_WIRE_24,
		 clr => SYNTHESIZED_WIRE_59,
		 Q => GDFX_TEMP_SIGNAL_3);


SYNTHESIZED_WIRE_59 <= CLK_50MHz OR SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_23 <= Q31 AND Q22;


b2v_inst39 : edgeing
PORT MAP(clk => CLK_50MHz,
		 D_in => SYNTHESIZED_WIRE_27,
		 Q => SYNTHESIZED_WIRE_18);


b2v_inst40 : edgeing
PORT MAP(clk => CLK_50MHz,
		 D_in => SYNTHESIZED_WIRE_56,
		 Q => SYNTHESIZED_WIRE_10);


b2v_inst41 : edgeing
PORT MAP(clk => CLK_50MHz,
		 D_in => SYNTHESIZED_WIRE_29,
		 Q => SYNTHESIZED_WIRE_19);


b2v_inst468 : bcd_to_7seg
PORT MAP(BCD_in => GDFX_TEMP_SIGNAL_4,
		 Seg_out => SYNTHESIZED_WIRE_60);


b2v_inst469 : bcd_to_7seg
PORT MAP(BCD_in => GDFX_TEMP_SIGNAL_5,
		 Seg_out => SYNTHESIZED_WIRE_61);


b2v_inst470 : bcd_to_7seg
PORT MAP(BCD_in => GDFX_TEMP_SIGNAL_6,
		 Seg_out => SYNTHESIZED_WIRE_62);


b2v_inst471 : bcd_to_7seg
PORT MAP(BCD_in => GDFX_TEMP_SIGNAL_7,
		 Seg_out => SYNTHESIZED_WIRE_63);


Q0 <= GDFX_TEMP_SIGNAL_0(0);
Q1 <= GDFX_TEMP_SIGNAL_0(1);
Q10 <= GDFX_TEMP_SIGNAL_1(0);
Q11 <= GDFX_TEMP_SIGNAL_1(1);
Q12 <= GDFX_TEMP_SIGNAL_1(2);
Q13 <= GDFX_TEMP_SIGNAL_1(3);
Q2 <= GDFX_TEMP_SIGNAL_0(2);
Q20 <= GDFX_TEMP_SIGNAL_2(0);
Q21 <= GDFX_TEMP_SIGNAL_2(1);
Q22 <= GDFX_TEMP_SIGNAL_2(2);
Q23 <= GDFX_TEMP_SIGNAL_2(3);
Q3 <= GDFX_TEMP_SIGNAL_0(3);
Q30 <= GDFX_TEMP_SIGNAL_3(0);
Q31 <= GDFX_TEMP_SIGNAL_3(1);
Q32 <= GDFX_TEMP_SIGNAL_3(2);
Q33 <= GDFX_TEMP_SIGNAL_3(3);
END bdf_type;